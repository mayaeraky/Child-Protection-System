LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SWITCHING IS PORT(
SWITCH1:IN STD_LOGIC;
OUTPUT1:OUT STD_LOGIC);
END SWITCHING;


ARCHITECTURE FUNCTION1 OF SWITCHING IS
BEGIN
WITH SWITCH1 SELECT
OUTPUT1<= '1' WHEN '1',
			 '0' WHEN OTHERS;
END FUNCTION1;